LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY vector_memory IS
	PORT (
		
		);
END vector_memory;

ARCHITECTURE comportamento OF vector_memory IS

BEGIN


END comportamento;