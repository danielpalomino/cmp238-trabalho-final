LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY difference IS
	PORT (
		
		);
END difference;

ARCHITECTURE comportamento OF difference IS

BEGIN


END comportamento;