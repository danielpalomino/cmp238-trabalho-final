LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE VECTOR_LIBRARY IS
	
	TYPE vector IS ARRAY (0 TO 1) OF STD_LOGIC_VECTOR(7 DOWNTO 0);	

END VECTOR_LIBRARY;