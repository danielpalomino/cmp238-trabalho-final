LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE VECTOR_LIBRARY IS

	TYPE motion_vector IS ARRAY (0 TO 1) OF STD_LOGIC_VECTOR(7 DOWNTO 0);

	COMPONENT mediana IS
		PORT (
			a, b, c : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			s : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		);
	END COMPONENT;


END VECTOR_LIBRARY;
