LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY comparator IS
	PORT (
		
		);
END comparator;

ARCHITECTURE comportamento OF comparator IS

BEGIN


END comportamento;