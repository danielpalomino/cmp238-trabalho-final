LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY vector_predictor IS
	PORT (
		
		);
END vector_predictor;

ARCHITECTURE comportamento OF vector_predictor IS

BEGIN


END comportamento;